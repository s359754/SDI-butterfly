
library IEEE;
use IEEE.std_logic_1164.all; --  libreria IEEE con definizione tipi standard logic
use IEEE.numeric_std.all;


entity BFLY_TOP_ENTITY is
port( 

);
end	BFLY_TOP_ENTITY;

---------------------------------------------

architecture structural of BFLY_TOP_ENTITY is
	
	component 
	
	
	begin
	
end structural;
 
